15 15 23 27 8 
W 12 11 9 5 23 
R 12 0 11 4 23 
R 14 1 11 4 23 
O 5 7 7 4 23 
R 13 7 11 4 23 
R 14 0 11 4 23 
O 0 8 4 4 23 
O 1 5 7 4 23 
O 9 10 4 4 23 
O 4 4 4 4 23 
A 6 7 4 4 23 
R 14 3 11 4 23 
A 0 14 4 4 23 
S 7 3 5 4 7 
R 9 0 11 4 3 
Z 10 6 2 1 23 
X 8 5 99 0 23 
T 14 8 0 0 23 
X 2 4 99 0 23 
G 3 7 0 0 23 
X 10 10 99 0 23 
T 3 8 0 0 23 
X 9 11 99 0 15 
X 1 0 99 0 12 
G 2 6 0 0 7 
X 7 10 99 0 7 
X 0 0 99 0 0 
#ZAPIS GRY WIRTUALNY SWIAT v3.0#
#Damian Jankowski s188597#
#znak polX polY sila inicjatywa wiek#
#[A]ntylopa [C]zlowiek [S]uperman [L]is [O]wca [W]ilk [Z]olw#
#[B]arszcz [G]uarana [M]lecz [T]rawa [X]Wilczejagody [R]CyberOwca#
#Superman - czlowiek z wlaczona umiejetnoscia#
